Howard Jones@HOWARDJONES-PC.3040:1444140520