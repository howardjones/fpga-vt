
constant BITS_PER_COLOUR : integer := 2;
constant CHAR_PER_LINE : integer := 80;
constant LINES_PER_SCREEN : integer := 25;

